LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY le_shift_entity IS
  PORT (
  );
END le_shift_entity;

ARCHITECTURE le_shift_architecture OF le_shift_entity IS
BEGIN
END le_shift_entity;