LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY boilerplate_entity IS
	PORT (
	);
END boilerplate_entity;

ARCHITECTURE boilerplate_architecture OF boilerplate_entity IS
BEGIN
END boilerplate_architecture;